module transmitter (
  input clk100_i,
  input rstn_i,
  input start,
  input data,
  output busy,
  output tx
);

endmodule
